/****************************************************************
/*
/*  Description:
/*              main FSM control of huffman coding process
/*  Author:
/*              Guozhu Xin
/*  Date:
/*              2017/7/11
/*  Email:
/*              spikexin@outlook.com
******************************************************************/

module HuffmanCode (
  input       clk,
  
  )
